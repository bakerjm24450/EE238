// Model of the Thunderbird turn signal.
// Turn-signal follows a simple pattern
module turnSignal(input logic clk,
                  input logic reset,
                  input logic signal,
                  output logic sa,
                  output logic sb,
                  output logic sc);
  

endmodule
