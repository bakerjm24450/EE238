// Seven-segment driver. Outputs hex values
module sevenSegDriver(input logic [3:0] digit,
			output logic ca,
			output logic cb,
			output logic cc,
			output logic cd,
			output logic ce,
			output logic cf,
			output logic cg);

	// FIXME -- Add your implementation here
	
endmodule
